library verilog;
use verilog.vl_types.all;
entity TM is
    generic(
        t               : integer := 1
    );
end TM;
