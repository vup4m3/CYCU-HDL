module Spi_Ctrl(
  input spi_en,
  input spi_clk,
  input [23:0]spi_wdata,
  input aluop_st,
  input rst
    
);


endmodule // Spi_Ctrl